

module fifo#(parameter WIDTH = 22 , parameter DEPTH=13)();

endmodule 