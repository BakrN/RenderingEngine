
module ren_top(); 

endmodule 