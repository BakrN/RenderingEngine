module ren_cu (
) ; 
    



  
endmodule 