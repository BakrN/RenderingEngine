`include "ren_defines.svh"

module ren_raster_queue( 
    // fifo info 
    i_write ,  
    i_tile , 
    o_tile ,  
); 
    input logic i_write, 
    input tile_t i_tile ; 
    input tile_t o_tile ; 
    


endmodule; 