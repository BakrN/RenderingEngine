module ren_cu (
    clk, 
    i_en ,  
    i_cmd , 
    // info 
    o_ack , 
) ; 
    



  
endmodule 